library verilog;
use verilog.vl_types.all;
entity Layer1_sv_unit is
end Layer1_sv_unit;
