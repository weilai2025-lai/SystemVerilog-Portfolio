library verilog;
use verilog.vl_types.all;
entity nn_config_pkg is
end nn_config_pkg;
