library verilog;
use verilog.vl_types.all;
entity neuron_opt_sv_unit is
end neuron_opt_sv_unit;
