library verilog;
use verilog.vl_types.all;
entity altlvds_rx is
    generic(
        number_of_channels: integer := 1;
        deserialization_factor: integer := 4;
        registered_output: string  := "ON";
        inclock_period  : integer := 10000;
        inclock_boost   : vl_notype;
        cds_mode        : string  := "UNUSED";
        intended_device_family: string  := "Stratix";
        input_data_rate : integer := 0;
        inclock_data_alignment: string  := "UNUSED";
        registered_data_align_input: string  := "ON";
        common_rx_tx_pll: string  := "ON";
        enable_dpa_mode : string  := "OFF";
        enable_dpa_calibration: string  := "ON";
        enable_dpa_pll_calibration: string  := "OFF";
        enable_dpa_fifo : string  := "ON";
        use_dpll_rawperror: string  := "OFF";
        use_coreclock_input: string  := "OFF";
        dpll_lock_count : integer := 0;
        dpll_lock_window: integer := 0;
        outclock_resource: string  := "AUTO";
        data_align_rollover: vl_notype;
        lose_lock_on_one_change: string  := "OFF";
        reset_fifo_at_first_lock: string  := "ON";
        use_external_pll: string  := "OFF";
        implement_in_les: string  := "OFF";
        buffer_implementation: string  := "RAM";
        port_rx_data_align: string  := "PORT_CONNECTIVITY";
        port_rx_channel_data_align: string  := "PORT_CONNECTIVITY";
        pll_operation_mode: string  := "NORMAL";
        x_on_bitslip    : string  := "ON";
        use_no_phase_shift: string  := "ON";
        rx_align_data_reg: string  := "RISING_EDGE";
        inclock_phase_shift: integer := 0;
        enable_soft_cdr_mode: string  := "OFF";
        sim_dpa_output_clock_phase_shift: integer := 0;
        sim_dpa_is_negative_ppm_drift: string  := "OFF";
        sim_dpa_net_ppm_variation: integer := 0;
        enable_dpa_align_to_rising_edge_only: string  := "OFF";
        enable_dpa_initial_phase_selection: string  := "OFF";
        dpa_initial_phase_value: integer := 0;
        pll_self_reset_on_loss_lock: string  := "OFF";
        refclk_frequency: string  := "UNUSED";
        enable_clock_pin_mode: string  := "UNUSED";
        data_rate       : string  := "UNUSED";
        lpm_hint        : string  := "UNUSED";
        lpm_type        : string  := "altlvds_rx";
        lvds_rx_reg_setting: string  := "ON";
        clk_src_is_pll  : string  := "off";
        STRATIX_RX_STYLE: vl_notype;
        STRATIXGX_DPA_RX_STYLE: vl_notype;
        STRATIXII_RX_STYLE: vl_notype;
        CYCLONE_RX_STYLE: vl_notype;
        CYCLONEII_RX_STYLE: vl_notype;
        STRATIXIII_RX_STYLE: vl_notype;
        ARRIAII_RX_STYLE: vl_notype;
        STRATIXV_RX_STYLE: vl_notype;
        CYCLONEIII_RX_STYLE: vl_notype;
        FAMILY_HAS_FLEXIBLE_LVDS: vl_notype;
        FAMILY_HAS_STRATIX_STYLE_PLL: vl_notype;
        FAMILY_HAS_STRATIXII_STYLE_PLL: vl_notype;
        FAMILY_HAS_STRATIXIII_STYLE_PLL: vl_notype;
        INT_CLOCK_BOOST : vl_notype;
        PLL_M_VALUE     : vl_notype;
        PLL_D_VALUE     : vl_notype;
        VSERIES_FAMILY  : vl_notype;
        STRATIX_INCLOCK_BOOST: vl_notype;
        PHASE_SHIFT     : vl_notype;
        STXII_PHASE_SHIFT: vl_notype;
        STXII_LE_PHASE_SHIFT: vl_notype;
        STXIII_LE_PHASE_SHIFT: vl_notype;
        REGISTER_WIDTH  : vl_notype;
        CLOCK_PERIOD    : vl_notype;
        FAST_CLK_ENA_PHASE_SHIFT: vl_notype;
        use_dpa_calibration: vl_notype
    );
    port(
        rx_in           : in     vl_logic_vector;
        rx_inclock      : in     vl_logic;
        rx_syncclock    : in     vl_logic;
        rx_dpaclock     : in     vl_logic;
        rx_readclock    : in     vl_logic;
        rx_enable       : in     vl_logic;
        rx_deskew       : in     vl_logic;
        rx_pll_enable   : in     vl_logic;
        rx_data_align   : in     vl_logic;
        rx_data_align_reset: in     vl_logic;
        rx_reset        : in     vl_logic_vector;
        rx_dpll_reset   : in     vl_logic_vector;
        rx_dpll_hold    : in     vl_logic_vector;
        rx_dpll_enable  : in     vl_logic_vector;
        rx_fifo_reset   : in     vl_logic_vector;
        rx_channel_data_align: in     vl_logic_vector;
        rx_cda_reset    : in     vl_logic_vector;
        rx_coreclk      : in     vl_logic_vector;
        pll_areset      : in     vl_logic;
        pll_phasedone   : in     vl_logic;
        dpa_pll_recal   : in     vl_logic;
        rx_dpa_lock_reset: in     vl_logic_vector;
        rx_out          : out    vl_logic_vector;
        rx_outclock     : out    vl_logic;
        rx_locked       : out    vl_logic;
        rx_dpa_locked   : out    vl_logic_vector;
        rx_cda_max      : out    vl_logic_vector;
        rx_divfwdclk    : out    vl_logic_vector;
        pll_phasestep   : out    vl_logic;
        pll_phaseupdown : out    vl_logic;
        pll_phasecounterselect: out    vl_logic_vector(3 downto 0);
        pll_scanclk     : out    vl_logic;
        dpa_pll_cal_busy: out    vl_logic;
        rx_data_reset   : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of number_of_channels : constant is 1;
    attribute mti_svvh_generic_type of deserialization_factor : constant is 1;
    attribute mti_svvh_generic_type of registered_output : constant is 1;
    attribute mti_svvh_generic_type of inclock_period : constant is 1;
    attribute mti_svvh_generic_type of inclock_boost : constant is 3;
    attribute mti_svvh_generic_type of cds_mode : constant is 1;
    attribute mti_svvh_generic_type of intended_device_family : constant is 1;
    attribute mti_svvh_generic_type of input_data_rate : constant is 1;
    attribute mti_svvh_generic_type of inclock_data_alignment : constant is 1;
    attribute mti_svvh_generic_type of registered_data_align_input : constant is 1;
    attribute mti_svvh_generic_type of common_rx_tx_pll : constant is 1;
    attribute mti_svvh_generic_type of enable_dpa_mode : constant is 1;
    attribute mti_svvh_generic_type of enable_dpa_calibration : constant is 1;
    attribute mti_svvh_generic_type of enable_dpa_pll_calibration : constant is 1;
    attribute mti_svvh_generic_type of enable_dpa_fifo : constant is 1;
    attribute mti_svvh_generic_type of use_dpll_rawperror : constant is 1;
    attribute mti_svvh_generic_type of use_coreclock_input : constant is 1;
    attribute mti_svvh_generic_type of dpll_lock_count : constant is 1;
    attribute mti_svvh_generic_type of dpll_lock_window : constant is 1;
    attribute mti_svvh_generic_type of outclock_resource : constant is 1;
    attribute mti_svvh_generic_type of data_align_rollover : constant is 3;
    attribute mti_svvh_generic_type of lose_lock_on_one_change : constant is 1;
    attribute mti_svvh_generic_type of reset_fifo_at_first_lock : constant is 1;
    attribute mti_svvh_generic_type of use_external_pll : constant is 1;
    attribute mti_svvh_generic_type of implement_in_les : constant is 1;
    attribute mti_svvh_generic_type of buffer_implementation : constant is 1;
    attribute mti_svvh_generic_type of port_rx_data_align : constant is 1;
    attribute mti_svvh_generic_type of port_rx_channel_data_align : constant is 1;
    attribute mti_svvh_generic_type of pll_operation_mode : constant is 1;
    attribute mti_svvh_generic_type of x_on_bitslip : constant is 1;
    attribute mti_svvh_generic_type of use_no_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of rx_align_data_reg : constant is 1;
    attribute mti_svvh_generic_type of inclock_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of enable_soft_cdr_mode : constant is 1;
    attribute mti_svvh_generic_type of sim_dpa_output_clock_phase_shift : constant is 1;
    attribute mti_svvh_generic_type of sim_dpa_is_negative_ppm_drift : constant is 1;
    attribute mti_svvh_generic_type of sim_dpa_net_ppm_variation : constant is 1;
    attribute mti_svvh_generic_type of enable_dpa_align_to_rising_edge_only : constant is 1;
    attribute mti_svvh_generic_type of enable_dpa_initial_phase_selection : constant is 1;
    attribute mti_svvh_generic_type of dpa_initial_phase_value : constant is 1;
    attribute mti_svvh_generic_type of pll_self_reset_on_loss_lock : constant is 1;
    attribute mti_svvh_generic_type of refclk_frequency : constant is 1;
    attribute mti_svvh_generic_type of enable_clock_pin_mode : constant is 1;
    attribute mti_svvh_generic_type of data_rate : constant is 1;
    attribute mti_svvh_generic_type of lpm_hint : constant is 1;
    attribute mti_svvh_generic_type of lpm_type : constant is 1;
    attribute mti_svvh_generic_type of lvds_rx_reg_setting : constant is 1;
    attribute mti_svvh_generic_type of clk_src_is_pll : constant is 1;
    attribute mti_svvh_generic_type of STRATIX_RX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of STRATIXGX_DPA_RX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of STRATIXII_RX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of CYCLONE_RX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of CYCLONEII_RX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of STRATIXIII_RX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of ARRIAII_RX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of STRATIXV_RX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of CYCLONEIII_RX_STYLE : constant is 3;
    attribute mti_svvh_generic_type of FAMILY_HAS_FLEXIBLE_LVDS : constant is 3;
    attribute mti_svvh_generic_type of FAMILY_HAS_STRATIX_STYLE_PLL : constant is 3;
    attribute mti_svvh_generic_type of FAMILY_HAS_STRATIXII_STYLE_PLL : constant is 3;
    attribute mti_svvh_generic_type of FAMILY_HAS_STRATIXIII_STYLE_PLL : constant is 3;
    attribute mti_svvh_generic_type of INT_CLOCK_BOOST : constant is 3;
    attribute mti_svvh_generic_type of PLL_M_VALUE : constant is 3;
    attribute mti_svvh_generic_type of PLL_D_VALUE : constant is 3;
    attribute mti_svvh_generic_type of VSERIES_FAMILY : constant is 3;
    attribute mti_svvh_generic_type of STRATIX_INCLOCK_BOOST : constant is 3;
    attribute mti_svvh_generic_type of PHASE_SHIFT : constant is 3;
    attribute mti_svvh_generic_type of STXII_PHASE_SHIFT : constant is 3;
    attribute mti_svvh_generic_type of STXII_LE_PHASE_SHIFT : constant is 3;
    attribute mti_svvh_generic_type of STXIII_LE_PHASE_SHIFT : constant is 3;
    attribute mti_svvh_generic_type of REGISTER_WIDTH : constant is 3;
    attribute mti_svvh_generic_type of CLOCK_PERIOD : constant is 3;
    attribute mti_svvh_generic_type of FAST_CLK_ENA_PHASE_SHIFT : constant is 3;
    attribute mti_svvh_generic_type of use_dpa_calibration : constant is 3;
end altlvds_rx;
