library verilog;
use verilog.vl_types.all;
entity Layer2_sv_unit is
end Layer2_sv_unit;
