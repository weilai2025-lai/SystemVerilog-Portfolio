library verilog;
use verilog.vl_types.all;
entity tb_neuron_opt_sv_unit is
end tb_neuron_opt_sv_unit;
