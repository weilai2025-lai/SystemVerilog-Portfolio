library verilog;
use verilog.vl_types.all;
entity Layer3_sv_unit is
end Layer3_sv_unit;
