library verilog;
use verilog.vl_types.all;
entity sig_rom_sv_unit is
end sig_rom_sv_unit;
