library verilog;
use verilog.vl_types.all;
entity dnn_sv_unit is
end dnn_sv_unit;
