library verilog;
use verilog.vl_types.all;
entity weight_memory_opt_sv_unit is
end weight_memory_opt_sv_unit;
