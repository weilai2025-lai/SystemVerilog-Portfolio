library verilog;
use verilog.vl_types.all;
entity weight_memory_sv_unit is
end weight_memory_sv_unit;
