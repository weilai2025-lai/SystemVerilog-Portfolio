library verilog;
use verilog.vl_types.all;
entity Layer4_sv_unit is
end Layer4_sv_unit;
