library verilog;
use verilog.vl_types.all;
entity tb_dnn_sv_unit is
end tb_dnn_sv_unit;
