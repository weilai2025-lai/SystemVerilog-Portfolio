library verilog;
use verilog.vl_types.all;
entity neuron_sv_unit is
end neuron_sv_unit;
