library verilog;
use verilog.vl_types.all;
entity maxfinder_sv_unit is
end maxfinder_sv_unit;
